library verilog;
use verilog.vl_types.all;
entity display_encoder_vlg_vec_tst is
end display_encoder_vlg_vec_tst;
