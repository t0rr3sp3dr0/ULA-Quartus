library verilog;
use verilog.vl_types.all;
entity placa_ULA_vlg_vec_tst is
end placa_ULA_vlg_vec_tst;
