library verilog;
use verilog.vl_types.all;
entity XOR30_vlg_vec_tst is
end XOR30_vlg_vec_tst;
