library verilog;
use verilog.vl_types.all;
entity BCD_demux_vlg_vec_tst is
end BCD_demux_vlg_vec_tst;
