library verilog;
use verilog.vl_types.all;
entity DEMUX_vlg_vec_tst is
end DEMUX_vlg_vec_tst;
