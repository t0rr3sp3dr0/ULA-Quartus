library verilog;
use verilog.vl_types.all;
entity b2d_vlg_check_tst is
    port(
        \_0000\         : in     vl_logic;
        \_1XXX\         : in     vl_logic;
        \_0001\         : in     vl_logic;
        \_0010\         : in     vl_logic;
        \_0011\         : in     vl_logic;
        \_0100\         : in     vl_logic;
        \_0101\         : in     vl_logic;
        \_0110\         : in     vl_logic;
        \_0111\         : in     vl_logic;
        \_1000\         : in     vl_logic;
        \_1001\         : in     vl_logic;
        \_1010\         : in     vl_logic;
        \_1011\         : in     vl_logic;
        \_1100\         : in     vl_logic;
        \_1101\         : in     vl_logic;
        \_1110\         : in     vl_logic;
        \_1111\         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end b2d_vlg_check_tst;
