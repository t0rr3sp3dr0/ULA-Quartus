library verilog;
use verilog.vl_types.all;
entity b2d_vlg_vec_tst is
end b2d_vlg_vec_tst;
