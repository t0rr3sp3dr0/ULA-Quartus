library verilog;
use verilog.vl_types.all;
entity inversor_vlg_vec_tst is
end inversor_vlg_vec_tst;
