library verilog;
use verilog.vl_types.all;
entity b2d is
    port(
        \_0000\         : out    vl_logic;
        E               : in     vl_logic_vector(3 downto 0);
        \_0001\         : out    vl_logic;
        \_0010\         : out    vl_logic;
        \_0011\         : out    vl_logic;
        \_0100\         : out    vl_logic;
        \_0101\         : out    vl_logic;
        \_0110\         : out    vl_logic;
        \_0111\         : out    vl_logic;
        \_1000\         : out    vl_logic;
        \_1001\         : out    vl_logic;
        \_1010\         : out    vl_logic;
        \_1011\         : out    vl_logic;
        \_1100\         : out    vl_logic;
        \_1101\         : out    vl_logic;
        \_1110\         : out    vl_logic;
        \_1111\         : out    vl_logic;
        \_1XXX\         : out    vl_logic
    );
end b2d;
