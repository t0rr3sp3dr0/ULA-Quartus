library verilog;
use verilog.vl_types.all;
entity AND30_vlg_vec_tst is
end AND30_vlg_vec_tst;
