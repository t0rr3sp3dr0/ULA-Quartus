library verilog;
use verilog.vl_types.all;
entity placa_BCD_vlg_vec_tst is
end placa_BCD_vlg_vec_tst;
