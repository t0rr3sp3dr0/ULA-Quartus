library verilog;
use verilog.vl_types.all;
entity BCD_demux is
    port(
        \_0\            : out    vl_logic;
        S               : in     vl_logic_vector(3 downto 0);
        \_1\            : out    vl_logic;
        \_2\            : out    vl_logic;
        \_3\            : out    vl_logic;
        \_4\            : out    vl_logic;
        \_5\            : out    vl_logic;
        \_6\            : out    vl_logic;
        \_7\            : out    vl_logic;
        \_8\            : out    vl_logic;
        \_9\            : out    vl_logic
    );
end BCD_demux;
