library verilog;
use verilog.vl_types.all;
entity BCD_demux_vlg_check_tst is
    port(
        \_0\            : in     vl_logic;
        \_1\            : in     vl_logic;
        \_2\            : in     vl_logic;
        \_3\            : in     vl_logic;
        \_4\            : in     vl_logic;
        \_5\            : in     vl_logic;
        \_6\            : in     vl_logic;
        \_7\            : in     vl_logic;
        \_8\            : in     vl_logic;
        \_9\            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end BCD_demux_vlg_check_tst;
