library verilog;
use verilog.vl_types.all;
entity display_encoder is
    port(
        display_a       : out    vl_logic;
        D               : in     vl_logic;
        \_4\            : in     vl_logic;
        \_1\            : in     vl_logic;
        B               : in     vl_logic;
        display_b       : out    vl_logic;
        F               : in     vl_logic;
        C               : in     vl_logic;
        E               : in     vl_logic;
        \_6\            : in     vl_logic;
        \_5\            : in     vl_logic;
        display_c       : out    vl_logic;
        \_2\            : in     vl_logic;
        display_d       : out    vl_logic;
        \_7\            : in     vl_logic;
        A               : in     vl_logic;
        display_e       : out    vl_logic;
        \_9\            : in     vl_logic;
        \_3\            : in     vl_logic;
        display_f       : out    vl_logic;
        display_g       : out    vl_logic;
        \_0\            : in     vl_logic;
        display_dp      : out    vl_logic;
        DP              : in     vl_logic;
        \_8\            : in     vl_logic
    );
end display_encoder;
