library verilog;
use verilog.vl_types.all;
entity display_encoder_vlg_sample_tst is
    port(
        \_0\            : in     vl_logic;
        \_1\            : in     vl_logic;
        \_2\            : in     vl_logic;
        \_3\            : in     vl_logic;
        \_4\            : in     vl_logic;
        \_5\            : in     vl_logic;
        \_6\            : in     vl_logic;
        \_7\            : in     vl_logic;
        \_8\            : in     vl_logic;
        \_9\            : in     vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        DP              : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end display_encoder_vlg_sample_tst;
