library verilog;
use verilog.vl_types.all;
entity BCD_decoder_vlg_vec_tst is
end BCD_decoder_vlg_vec_tst;
